program bathtub_test();
  
  task main();
    $info("Hello, world!");
  endtask : main
  
  initial main();
  
endprogram : bathtub_test